library verilog;
use verilog.vl_types.all;
entity compU8_vlg_vec_tst is
end compU8_vlg_vec_tst;
