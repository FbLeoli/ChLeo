library verilog;
use verilog.vl_types.all;
entity som_sub_sig_vlg_vec_tst is
end som_sub_sig_vlg_vec_tst;
