library verilog;
use verilog.vl_types.all;
entity micro_vlg_vec_tst is
end micro_vlg_vec_tst;
