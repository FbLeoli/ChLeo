library verilog;
use verilog.vl_types.all;
entity comp8_vlg_vec_tst is
end comp8_vlg_vec_tst;
